// ============================================================================
// lfsr32.sv
// 매 클럭마다 값이 한 칸씩 왼쪽으로 밀리고, 
// 맨 오른쪽에는 몇개 비트를 XOR한 값이 새로 들어옴 (XOR를 사용해야 0과 1이 골고루 섞긴 긴 주기 패턴이 나와 난수 사용 가능)
// 리셋이 0이면 정해둔 시작값으로 다시 시작함
//============================================================================
module lfsr32(
  input  logic clk,
  input  logic rst_n,
  output logic [31:0] q // 바깥으로 보여줄 32비트 현재 값
);
  logic [31:0] r; // 내부에서 값 들고 있는 32비트 레지스터

  // 클럭이 1로 올라갈 때 또는 리셋이 1->0으로 내려갈 때 반응 
  always_ff @(posedge clk or negedge rst_n) begin 
    if(!rst_n) r <= 32'h1ACE_B00C; // 리셋이 0이면, 시작값으로 설정
    else       r <= {r[30:0], r[31]^r[21]^r[1]^r[0]};
    // 리셋이 아니면 매 클럭마다, r을 한 칸 왼쪽으로 민 다음, 맨 오른쪽 비트에는 값들을 xor한 값을 넣음
    // 이렇게 패턴이 반복되면서 난수처럼 보이는 수열이 나옴
  end
  assign q = r; // 내부 값 r을 그대로 출력 q에 연결 
endmodule
